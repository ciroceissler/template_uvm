`ifndef TEMPLATE_TYPES_SVH
`define TEMPLATE_TYPES_SVH

typedef virtual template_if template_vif_t;

`endif // TEMPLATE_TYPES_SVH

