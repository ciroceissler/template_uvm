`infdef TEMPLATE_TYPES_SV

  typedef virtual template_if template_vif_t;

`endif // TEMPLATE_TYPES_SV
