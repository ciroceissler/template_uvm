`ifndef TEMPLATE_FUNCOV_SVH
`define TEMPLATE_FUNCOV_SVH

class template_funcov;
endclass : template_funcov

`endif // TEMPLATE_FUNCOV_SVH

