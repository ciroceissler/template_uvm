module template (
  input  clk,
  input  rst,
  input  data_i,
  output data_o
);

  assign data_o = data_i; 

endmodule : template

