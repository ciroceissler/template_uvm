module template_tb;

  // +--------------------------------------------------------------------------
  // | local variables
  // +--------------------------------------------------------------------------
  logic clk;
  logic rst;
  logic data_i;
  logic data_o;

  // +--------------------------------------------------------------------------
  // | instantiate modules
  // +--------------------------------------------------------------------------
  template uu_template (
    .clk    (clk),
    .rst    (rst),
    .data_i (data_i),
    .data_o (data_o)
  );

  // +--------------------------------------------------------------------------
  // | TASK: run_clk
  // +--------------------------------------------------------------------------
  task run_clk();
    forever begin
      #5 clk <= ~clk;
    end
  endtask : run_clk

  // +--------------------------------------------------------------------------
  // | TASK: run_reset
  // +--------------------------------------------------------------------------
  task run_reset();
    #10 rst = 1'b1;
    #10 rst = 1'b0;
  endtask : run_reset

  // +--------------------------------------------------------------------------
  // | TASK: run
  // +--------------------------------------------------------------------------
  task run(int unsigned num);
    for (int i = 0; i < num; i++) begin
      data_i <= $urandom;

      @(posedge clk);
    end
  endtask : run

  // +--------------------------------------------------------------------------
  // | BLOCK: main block
  // +--------------------------------------------------------------------------
  initial begin
    int unsigned num;

    clk    = '0;
    rst    = '0;
    data_i = '0;

    if (!$value$plusargs ("num=%d", num))
      num = 1000;

    fork
      run_clk();
      run_reset();
    join_none

    run(num);

    $finish;
  end

endmodule : template_tb

