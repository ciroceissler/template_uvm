package template_agent_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"
  
  `include "template_types.sv"
  `include "template_sqc_item.sv"
  `include "template_sqc_base.sv"
  `include "template_sqc_api.sv"
  `include "template_sequencer.sv"
  `include "template_driver.sv"
  `include "template_monitor.sv"
  `include "template_agent_config.sv"
  `include "template_agent.sv"

endpackage : template_agent_pkg;
