class template_funcov;
endclass : template_funcov
