`include "template_test_bypass.sv"
