`ifndef TEMPLATE_TEST_LIST_SVH
`define TEMPLATE_TEST_LIST_SVH

`include "template_report_server.svh"
`include "template_test_report.svh"
`include "template_test_base.svh"
`include "template_test_bypass.svh"

`endif // TEMPLATE_TEST_LIST_SVH

