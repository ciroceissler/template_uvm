module template (
  input  clk,
  input  rst,
  input  data_i,
  output data_o
);

  // NOTE(ciroceissler): stub

endmodule : template

