package template_agent_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "template_types.svh"
  `include "template_agent_config.svh"
  `include "template_sqc_item.svh"
  `include "template_sqc_base.svh"
  `include "template_sqc_api.svh"
  `include "template_sequencer.svh"
  `include "template_driver.svh"
  `include "template_monitor.svh"
  `include "template_agent.svh"

endpackage : template_agent_pkg

